`ifndef __DTM__
`define __DTM__

module DTM
(


);








endmodule


`endif