module multi(
ain,bin,ss,su,uu,cout,rstn,clk);

input ss,su,uu;
input[31:0] ain,bin;
output[31:0] cout;





endmodule
