`ifndef __DM__
`define __DM__

module DM
(


);







endmodule


`endif