`ifndef __TAP_CTRL__
`define __TAP_CTRL__

module TAP_ctrl
(
    input wire tck,//t-clk
    input wire trst,//t-reset
    input wire tms,//t-mode select

);









endmodule


`endif