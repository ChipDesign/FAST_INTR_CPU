`infdef __PARAMETERS__
`define __PARAMETERS__
    parameter INTR_SIZE = 128;
    parameter INTR_WIDTH =7;
    parameter INTR_SIZE_by32 =2;
`endif