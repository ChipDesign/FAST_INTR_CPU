module Pri_elem_8(
  input        clock,
  input        reset,
  output [4:0] io_pri,
  input  [4:0] io_pri_update,
  input        io_pri_update_sig
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] Pri; // @[Priority_agent.scala 21:18]
  assign io_pri = Pri; // @[Priority_agent.scala 31:9]
  always @(posedge clock) begin
    if (reset) begin // @[Priority_agent.scala 21:18]
      Pri <= 5'h2; // @[Priority_agent.scala 21:18]
    end else if (io_pri_update_sig) begin // @[Priority_agent.scala 40:3]
      Pri <= io_pri_update; // @[Priority_agent.scala 40:7]
    end else if (io_pri_update_sig) begin // @[Priority_agent.scala 27:3]
      Pri <= io_pri_update; // @[Priority_agent.scala 28:8]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  Pri = _RAND_0[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Pri_elem_9(
  input        clock,
  input        reset,
  output [4:0] io_pri,
  input  [4:0] io_pri_update,
  input        io_pri_update_sig
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] Pri; // @[Priority_agent.scala 21:18]
  assign io_pri = Pri; // @[Priority_agent.scala 31:9]
  always @(posedge clock) begin
    if (reset) begin // @[Priority_agent.scala 21:18]
      Pri <= 5'h2; // @[Priority_agent.scala 21:18]
    end else if (io_pri_update_sig) begin // @[Priority_agent.scala 40:3]
      Pri <= io_pri_update; // @[Priority_agent.scala 40:7]
    end else if (io_pri_update_sig) begin // @[Priority_agent.scala 27:3]
      Pri <= io_pri_update; // @[Priority_agent.scala 28:8]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  Pri = _RAND_0[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Pri_elem_10(
  input        clock,
  input        reset,
  output [4:0] io_pri,
  input  [4:0] io_pri_update,
  input        io_pri_update_sig
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] Pri; // @[Priority_agent.scala 21:18]
  assign io_pri = Pri; // @[Priority_agent.scala 31:9]
  always @(posedge clock) begin
    if (reset) begin // @[Priority_agent.scala 21:18]
      Pri <= 5'h2; // @[Priority_agent.scala 21:18]
    end else if (io_pri_update_sig) begin // @[Priority_agent.scala 40:3]
      Pri <= io_pri_update; // @[Priority_agent.scala 40:7]
    end else if (io_pri_update_sig) begin // @[Priority_agent.scala 27:3]
      Pri <= io_pri_update; // @[Priority_agent.scala 28:8]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  Pri = _RAND_0[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Pri_elem_11(
  input        clock,
  input        reset,
  output [4:0] io_pri,
  input  [4:0] io_pri_update,
  input        io_pri_update_sig
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] Pri; // @[Priority_agent.scala 21:18]
  assign io_pri = Pri; // @[Priority_agent.scala 31:9]
  always @(posedge clock) begin
    if (reset) begin // @[Priority_agent.scala 21:18]
      Pri <= 5'h2; // @[Priority_agent.scala 21:18]
    end else if (io_pri_update_sig) begin // @[Priority_agent.scala 40:3]
      Pri <= io_pri_update; // @[Priority_agent.scala 40:7]
    end else if (io_pri_update_sig) begin // @[Priority_agent.scala 27:3]
      Pri <= io_pri_update; // @[Priority_agent.scala 28:8]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  Pri = _RAND_0[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Pri_elem_12(
  input        clock,
  input        reset,
  output [4:0] io_pri,
  input  [4:0] io_pri_update,
  input        io_pri_update_sig
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] Pri; // @[Priority_agent.scala 21:18]
  assign io_pri = Pri; // @[Priority_agent.scala 31:9]
  always @(posedge clock) begin
    if (reset) begin // @[Priority_agent.scala 21:18]
      Pri <= 5'h2; // @[Priority_agent.scala 21:18]
    end else if (io_pri_update_sig) begin // @[Priority_agent.scala 40:3]
      Pri <= io_pri_update; // @[Priority_agent.scala 40:7]
    end else if (io_pri_update_sig) begin // @[Priority_agent.scala 27:3]
      Pri <= io_pri_update; // @[Priority_agent.scala 28:8]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  Pri = _RAND_0[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Pri_elem_13(
  input        clock,
  input        reset,
  output [4:0] io_pri,
  input  [4:0] io_pri_update,
  input        io_pri_update_sig
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] Pri; // @[Priority_agent.scala 21:18]
  assign io_pri = Pri; // @[Priority_agent.scala 31:9]
  always @(posedge clock) begin
    if (reset) begin // @[Priority_agent.scala 21:18]
      Pri <= 5'h2; // @[Priority_agent.scala 21:18]
    end else if (io_pri_update_sig) begin // @[Priority_agent.scala 40:3]
      Pri <= io_pri_update; // @[Priority_agent.scala 40:7]
    end else if (io_pri_update_sig) begin // @[Priority_agent.scala 27:3]
      Pri <= io_pri_update; // @[Priority_agent.scala 28:8]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  Pri = _RAND_0[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Pri_elem_14(
  input        clock,
  input        reset,
  output [4:0] io_pri,
  input  [4:0] io_pri_update,
  input        io_pri_update_sig
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] Pri; // @[Priority_agent.scala 21:18]
  assign io_pri = Pri; // @[Priority_agent.scala 31:9]
  always @(posedge clock) begin
    if (reset) begin // @[Priority_agent.scala 21:18]
      Pri <= 5'h2; // @[Priority_agent.scala 21:18]
    end else if (io_pri_update_sig) begin // @[Priority_agent.scala 40:3]
      Pri <= io_pri_update; // @[Priority_agent.scala 40:7]
    end else if (io_pri_update_sig) begin // @[Priority_agent.scala 27:3]
      Pri <= io_pri_update; // @[Priority_agent.scala 28:8]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  Pri = _RAND_0[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Pri_elem_15(
  input        clock,
  input        reset,
  output [4:0] io_pri,
  input  [4:0] io_pri_update,
  input        io_pri_update_sig
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] Pri; // @[Priority_agent.scala 21:18]
  assign io_pri = Pri; // @[Priority_agent.scala 31:9]
  always @(posedge clock) begin
    if (reset) begin // @[Priority_agent.scala 21:18]
      Pri <= 5'h2; // @[Priority_agent.scala 21:18]
    end else if (io_pri_update_sig) begin // @[Priority_agent.scala 40:3]
      Pri <= io_pri_update; // @[Priority_agent.scala 40:7]
    end else if (io_pri_update_sig) begin // @[Priority_agent.scala 27:3]
      Pri <= io_pri_update; // @[Priority_agent.scala 28:8]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  Pri = _RAND_0[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module By_ID_sel(
  output       io_sel_sig_0,
  output       io_sel_sig_1,
  output       io_sel_sig_2,
  output       io_sel_sig_3,
  output       io_sel_sig_4,
  output       io_sel_sig_5,
  output       io_sel_sig_6,
  output       io_sel_sig_7,
  input  [3:0] io_ID_in
);
  assign io_sel_sig_0 = io_ID_in == 4'h8; // @[By_ID_sel.scala 21:31]
  assign io_sel_sig_1 = io_ID_in == 4'h9; // @[By_ID_sel.scala 21:31]
  assign io_sel_sig_2 = io_ID_in == 4'ha; // @[By_ID_sel.scala 21:31]
  assign io_sel_sig_3 = io_ID_in == 4'hb; // @[By_ID_sel.scala 21:31]
  assign io_sel_sig_4 = io_ID_in == 4'hc; // @[By_ID_sel.scala 21:31]
  assign io_sel_sig_5 = io_ID_in == 4'hd; // @[By_ID_sel.scala 21:31]
  assign io_sel_sig_6 = io_ID_in == 4'he; // @[By_ID_sel.scala 21:31]
  assign io_sel_sig_7 = io_ID_in == 4'hf; // @[By_ID_sel.scala 21:31]
endmodule
module Priority_agent(
  input        clock,
  input        reset,
  input        io_dyn_int_claim_sig,
  output [4:0] io_int_pri_0,
  output [4:0] io_int_pri_1,
  output [4:0] io_int_pri_2,
  output [4:0] io_int_pri_3,
  output [4:0] io_int_pri_4,
  output [4:0] io_int_pri_5,
  output [4:0] io_int_pri_6,
  output [4:0] io_int_pri_7,
  output [4:0] io_int_pri_8,
  output [4:0] io_int_pri_9,
  output [4:0] io_int_pri_10,
  output [4:0] io_int_pri_11,
  output [4:0] io_int_pri_12,
  output [4:0] io_int_pri_13,
  output [4:0] io_int_pri_14,
  output [4:0] io_int_pri_15,
  input        io_dyn_int_occ_sig,
  input  [3:0] io_dyn_int_occ_ID,
  input  [3:0] io_dyn_int_claim_ID
);
  wire  Pri_elem_8_clock; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_8_reset; // @[Priority_agent.scala 54:24]
  wire [4:0] Pri_elem_8_io_pri; // @[Priority_agent.scala 54:24]
  wire [4:0] Pri_elem_8_io_pri_update; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_8_io_pri_update_sig; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_9_clock; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_9_reset; // @[Priority_agent.scala 54:24]
  wire [4:0] Pri_elem_9_io_pri; // @[Priority_agent.scala 54:24]
  wire [4:0] Pri_elem_9_io_pri_update; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_9_io_pri_update_sig; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_10_clock; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_10_reset; // @[Priority_agent.scala 54:24]
  wire [4:0] Pri_elem_10_io_pri; // @[Priority_agent.scala 54:24]
  wire [4:0] Pri_elem_10_io_pri_update; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_10_io_pri_update_sig; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_11_clock; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_11_reset; // @[Priority_agent.scala 54:24]
  wire [4:0] Pri_elem_11_io_pri; // @[Priority_agent.scala 54:24]
  wire [4:0] Pri_elem_11_io_pri_update; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_11_io_pri_update_sig; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_12_clock; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_12_reset; // @[Priority_agent.scala 54:24]
  wire [4:0] Pri_elem_12_io_pri; // @[Priority_agent.scala 54:24]
  wire [4:0] Pri_elem_12_io_pri_update; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_12_io_pri_update_sig; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_13_clock; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_13_reset; // @[Priority_agent.scala 54:24]
  wire [4:0] Pri_elem_13_io_pri; // @[Priority_agent.scala 54:24]
  wire [4:0] Pri_elem_13_io_pri_update; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_13_io_pri_update_sig; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_14_clock; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_14_reset; // @[Priority_agent.scala 54:24]
  wire [4:0] Pri_elem_14_io_pri; // @[Priority_agent.scala 54:24]
  wire [4:0] Pri_elem_14_io_pri_update; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_14_io_pri_update_sig; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_15_clock; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_15_reset; // @[Priority_agent.scala 54:24]
  wire [4:0] Pri_elem_15_io_pri; // @[Priority_agent.scala 54:24]
  wire [4:0] Pri_elem_15_io_pri_update; // @[Priority_agent.scala 54:24]
  wire  Pri_elem_15_io_pri_update_sig; // @[Priority_agent.scala 54:24]
  wire  IntClaimSel_io_sel_sig_0; // @[Priority_agent.scala 59:25]
  wire  IntClaimSel_io_sel_sig_1; // @[Priority_agent.scala 59:25]
  wire  IntClaimSel_io_sel_sig_2; // @[Priority_agent.scala 59:25]
  wire  IntClaimSel_io_sel_sig_3; // @[Priority_agent.scala 59:25]
  wire  IntClaimSel_io_sel_sig_4; // @[Priority_agent.scala 59:25]
  wire  IntClaimSel_io_sel_sig_5; // @[Priority_agent.scala 59:25]
  wire  IntClaimSel_io_sel_sig_6; // @[Priority_agent.scala 59:25]
  wire  IntClaimSel_io_sel_sig_7; // @[Priority_agent.scala 59:25]
  wire [3:0] IntClaimSel_io_ID_in; // @[Priority_agent.scala 59:25]
  wire  IntOccSel_io_sel_sig_0; // @[Priority_agent.scala 60:23]
  wire  IntOccSel_io_sel_sig_1; // @[Priority_agent.scala 60:23]
  wire  IntOccSel_io_sel_sig_2; // @[Priority_agent.scala 60:23]
  wire  IntOccSel_io_sel_sig_3; // @[Priority_agent.scala 60:23]
  wire  IntOccSel_io_sel_sig_4; // @[Priority_agent.scala 60:23]
  wire  IntOccSel_io_sel_sig_5; // @[Priority_agent.scala 60:23]
  wire  IntOccSel_io_sel_sig_6; // @[Priority_agent.scala 60:23]
  wire  IntOccSel_io_sel_sig_7; // @[Priority_agent.scala 60:23]
  wire [3:0] IntOccSel_io_ID_in; // @[Priority_agent.scala 60:23]
  wire [4:0] _T_1 = IntOccSel_io_sel_sig_0 ? 5'h1f : 5'h0; // @[Bitwise.scala 77:12]
  wire [4:0] _T_2 = _T_1 & 5'h2; // @[Priority_agent.scala 94:73]
  wire  _T_4 = ~IntOccSel_io_sel_sig_0 & io_dyn_int_occ_sig; // @[Priority_agent.scala 95:50]
  wire [4:0] _T_6 = _T_4 ? 5'h1f : 5'h0; // @[Bitwise.scala 77:12]
  wire [4:0] DynamPriUpdate_0 = Pri_elem_8_io_pri + 5'h1; // @[Priority_agent.scala 103:44]
  wire [4:0] _T_7 = _T_6 & DynamPriUpdate_0; // @[Priority_agent.scala 95:64]
  wire [4:0] _T_12 = IntOccSel_io_sel_sig_1 ? 5'h1f : 5'h0; // @[Bitwise.scala 77:12]
  wire [4:0] _T_13 = _T_12 & 5'h2; // @[Priority_agent.scala 94:73]
  wire  _T_15 = ~IntOccSel_io_sel_sig_1 & io_dyn_int_occ_sig; // @[Priority_agent.scala 95:50]
  wire [4:0] _T_17 = _T_15 ? 5'h1f : 5'h0; // @[Bitwise.scala 77:12]
  wire [4:0] DynamPriUpdate_1 = Pri_elem_9_io_pri + 5'h1; // @[Priority_agent.scala 103:44]
  wire [4:0] _T_18 = _T_17 & DynamPriUpdate_1; // @[Priority_agent.scala 95:64]
  wire [4:0] _T_23 = IntOccSel_io_sel_sig_2 ? 5'h1f : 5'h0; // @[Bitwise.scala 77:12]
  wire [4:0] _T_24 = _T_23 & 5'h2; // @[Priority_agent.scala 94:73]
  wire  _T_26 = ~IntOccSel_io_sel_sig_2 & io_dyn_int_occ_sig; // @[Priority_agent.scala 95:50]
  wire [4:0] _T_28 = _T_26 ? 5'h1f : 5'h0; // @[Bitwise.scala 77:12]
  wire [4:0] DynamPriUpdate_2 = Pri_elem_10_io_pri + 5'h1; // @[Priority_agent.scala 103:44]
  wire [4:0] _T_29 = _T_28 & DynamPriUpdate_2; // @[Priority_agent.scala 95:64]
  wire [4:0] _T_34 = IntOccSel_io_sel_sig_3 ? 5'h1f : 5'h0; // @[Bitwise.scala 77:12]
  wire [4:0] _T_35 = _T_34 & 5'h2; // @[Priority_agent.scala 94:73]
  wire  _T_37 = ~IntOccSel_io_sel_sig_3 & io_dyn_int_occ_sig; // @[Priority_agent.scala 95:50]
  wire [4:0] _T_39 = _T_37 ? 5'h1f : 5'h0; // @[Bitwise.scala 77:12]
  wire [4:0] DynamPriUpdate_3 = Pri_elem_11_io_pri + 5'h1; // @[Priority_agent.scala 103:44]
  wire [4:0] _T_40 = _T_39 & DynamPriUpdate_3; // @[Priority_agent.scala 95:64]
  wire [4:0] _T_45 = IntOccSel_io_sel_sig_4 ? 5'h1f : 5'h0; // @[Bitwise.scala 77:12]
  wire [4:0] _T_46 = _T_45 & 5'h2; // @[Priority_agent.scala 94:73]
  wire  _T_48 = ~IntOccSel_io_sel_sig_4 & io_dyn_int_occ_sig; // @[Priority_agent.scala 95:50]
  wire [4:0] _T_50 = _T_48 ? 5'h1f : 5'h0; // @[Bitwise.scala 77:12]
  wire [4:0] DynamPriUpdate_4 = Pri_elem_12_io_pri + 5'h1; // @[Priority_agent.scala 103:44]
  wire [4:0] _T_51 = _T_50 & DynamPriUpdate_4; // @[Priority_agent.scala 95:64]
  wire [4:0] _T_56 = IntOccSel_io_sel_sig_5 ? 5'h1f : 5'h0; // @[Bitwise.scala 77:12]
  wire [4:0] _T_57 = _T_56 & 5'h2; // @[Priority_agent.scala 94:73]
  wire  _T_59 = ~IntOccSel_io_sel_sig_5 & io_dyn_int_occ_sig; // @[Priority_agent.scala 95:50]
  wire [4:0] _T_61 = _T_59 ? 5'h1f : 5'h0; // @[Bitwise.scala 77:12]
  wire [4:0] DynamPriUpdate_5 = Pri_elem_13_io_pri + 5'h1; // @[Priority_agent.scala 103:44]
  wire [4:0] _T_62 = _T_61 & DynamPriUpdate_5; // @[Priority_agent.scala 95:64]
  wire [4:0] _T_67 = IntOccSel_io_sel_sig_6 ? 5'h1f : 5'h0; // @[Bitwise.scala 77:12]
  wire [4:0] _T_68 = _T_67 & 5'h2; // @[Priority_agent.scala 94:73]
  wire  _T_70 = ~IntOccSel_io_sel_sig_6 & io_dyn_int_occ_sig; // @[Priority_agent.scala 95:50]
  wire [4:0] _T_72 = _T_70 ? 5'h1f : 5'h0; // @[Bitwise.scala 77:12]
  wire [4:0] DynamPriUpdate_6 = Pri_elem_14_io_pri + 5'h1; // @[Priority_agent.scala 103:44]
  wire [4:0] _T_73 = _T_72 & DynamPriUpdate_6; // @[Priority_agent.scala 95:64]
  wire [4:0] _T_78 = IntOccSel_io_sel_sig_7 ? 5'h1f : 5'h0; // @[Bitwise.scala 77:12]
  wire [4:0] _T_79 = _T_78 & 5'h2; // @[Priority_agent.scala 94:73]
  wire  _T_81 = ~IntOccSel_io_sel_sig_7 & io_dyn_int_occ_sig; // @[Priority_agent.scala 95:50]
  wire [4:0] _T_83 = _T_81 ? 5'h1f : 5'h0; // @[Bitwise.scala 77:12]
  wire [4:0] DynamPriUpdate_7 = Pri_elem_15_io_pri + 5'h1; // @[Priority_agent.scala 103:44]
  wire [4:0] _T_84 = _T_83 & DynamPriUpdate_7; // @[Priority_agent.scala 95:64]
  Pri_elem_8 Pri_elem_8 ( // @[Priority_agent.scala 54:24]
    .clock(Pri_elem_8_clock),
    .reset(Pri_elem_8_reset),
    .io_pri(Pri_elem_8_io_pri),
    .io_pri_update(Pri_elem_8_io_pri_update),
    .io_pri_update_sig(Pri_elem_8_io_pri_update_sig)
  );
  Pri_elem_9 Pri_elem_9 ( // @[Priority_agent.scala 54:24]
    .clock(Pri_elem_9_clock),
    .reset(Pri_elem_9_reset),
    .io_pri(Pri_elem_9_io_pri),
    .io_pri_update(Pri_elem_9_io_pri_update),
    .io_pri_update_sig(Pri_elem_9_io_pri_update_sig)
  );
  Pri_elem_10 Pri_elem_10 ( // @[Priority_agent.scala 54:24]
    .clock(Pri_elem_10_clock),
    .reset(Pri_elem_10_reset),
    .io_pri(Pri_elem_10_io_pri),
    .io_pri_update(Pri_elem_10_io_pri_update),
    .io_pri_update_sig(Pri_elem_10_io_pri_update_sig)
  );
  Pri_elem_11 Pri_elem_11 ( // @[Priority_agent.scala 54:24]
    .clock(Pri_elem_11_clock),
    .reset(Pri_elem_11_reset),
    .io_pri(Pri_elem_11_io_pri),
    .io_pri_update(Pri_elem_11_io_pri_update),
    .io_pri_update_sig(Pri_elem_11_io_pri_update_sig)
  );
  Pri_elem_12 Pri_elem_12 ( // @[Priority_agent.scala 54:24]
    .clock(Pri_elem_12_clock),
    .reset(Pri_elem_12_reset),
    .io_pri(Pri_elem_12_io_pri),
    .io_pri_update(Pri_elem_12_io_pri_update),
    .io_pri_update_sig(Pri_elem_12_io_pri_update_sig)
  );
  Pri_elem_13 Pri_elem_13 ( // @[Priority_agent.scala 54:24]
    .clock(Pri_elem_13_clock),
    .reset(Pri_elem_13_reset),
    .io_pri(Pri_elem_13_io_pri),
    .io_pri_update(Pri_elem_13_io_pri_update),
    .io_pri_update_sig(Pri_elem_13_io_pri_update_sig)
  );
  Pri_elem_14 Pri_elem_14 ( // @[Priority_agent.scala 54:24]
    .clock(Pri_elem_14_clock),
    .reset(Pri_elem_14_reset),
    .io_pri(Pri_elem_14_io_pri),
    .io_pri_update(Pri_elem_14_io_pri_update),
    .io_pri_update_sig(Pri_elem_14_io_pri_update_sig)
  );
  Pri_elem_15 Pri_elem_15 ( // @[Priority_agent.scala 54:24]
    .clock(Pri_elem_15_clock),
    .reset(Pri_elem_15_reset),
    .io_pri(Pri_elem_15_io_pri),
    .io_pri_update(Pri_elem_15_io_pri_update),
    .io_pri_update_sig(Pri_elem_15_io_pri_update_sig)
  );
  By_ID_sel IntClaimSel ( // @[Priority_agent.scala 59:25]
    .io_sel_sig_0(IntClaimSel_io_sel_sig_0),
    .io_sel_sig_1(IntClaimSel_io_sel_sig_1),
    .io_sel_sig_2(IntClaimSel_io_sel_sig_2),
    .io_sel_sig_3(IntClaimSel_io_sel_sig_3),
    .io_sel_sig_4(IntClaimSel_io_sel_sig_4),
    .io_sel_sig_5(IntClaimSel_io_sel_sig_5),
    .io_sel_sig_6(IntClaimSel_io_sel_sig_6),
    .io_sel_sig_7(IntClaimSel_io_sel_sig_7),
    .io_ID_in(IntClaimSel_io_ID_in)
  );
  By_ID_sel IntOccSel ( // @[Priority_agent.scala 60:23]
    .io_sel_sig_0(IntOccSel_io_sel_sig_0),
    .io_sel_sig_1(IntOccSel_io_sel_sig_1),
    .io_sel_sig_2(IntOccSel_io_sel_sig_2),
    .io_sel_sig_3(IntOccSel_io_sel_sig_3),
    .io_sel_sig_4(IntOccSel_io_sel_sig_4),
    .io_sel_sig_5(IntOccSel_io_sel_sig_5),
    .io_sel_sig_6(IntOccSel_io_sel_sig_6),
    .io_sel_sig_7(IntOccSel_io_sel_sig_7),
    .io_ID_in(IntOccSel_io_ID_in)
  );
  assign io_int_pri_0 = 5'h1; // @[Priority_agent.scala 75:18]
  assign io_int_pri_1 = 5'h1; // @[Priority_agent.scala 75:18]
  assign io_int_pri_2 = 5'h1; // @[Priority_agent.scala 75:18]
  assign io_int_pri_3 = 5'h1; // @[Priority_agent.scala 75:18]
  assign io_int_pri_4 = 5'h1; // @[Priority_agent.scala 75:18]
  assign io_int_pri_5 = 5'h1; // @[Priority_agent.scala 75:18]
  assign io_int_pri_6 = 5'h1; // @[Priority_agent.scala 75:18]
  assign io_int_pri_7 = 5'h1; // @[Priority_agent.scala 75:18]
  assign io_int_pri_8 = Pri_elem_8_io_pri; // @[Priority_agent.scala 78:31]
  assign io_int_pri_9 = Pri_elem_9_io_pri; // @[Priority_agent.scala 78:31]
  assign io_int_pri_10 = Pri_elem_10_io_pri; // @[Priority_agent.scala 78:31]
  assign io_int_pri_11 = Pri_elem_11_io_pri; // @[Priority_agent.scala 78:31]
  assign io_int_pri_12 = Pri_elem_12_io_pri; // @[Priority_agent.scala 78:31]
  assign io_int_pri_13 = Pri_elem_13_io_pri; // @[Priority_agent.scala 78:31]
  assign io_int_pri_14 = Pri_elem_14_io_pri; // @[Priority_agent.scala 78:31]
  assign io_int_pri_15 = Pri_elem_15_io_pri; // @[Priority_agent.scala 78:31]
  assign Pri_elem_8_clock = clock;
  assign Pri_elem_8_reset = reset;
  assign Pri_elem_8_io_pri_update = _T_2 | _T_7; // @[Priority_agent.scala 94:84]
  assign Pri_elem_8_io_pri_update_sig = io_dyn_int_occ_sig; // @[Priority_agent.scala 100:35]
  assign Pri_elem_9_clock = clock;
  assign Pri_elem_9_reset = reset;
  assign Pri_elem_9_io_pri_update = _T_13 | _T_18; // @[Priority_agent.scala 94:84]
  assign Pri_elem_9_io_pri_update_sig = io_dyn_int_occ_sig; // @[Priority_agent.scala 100:35]
  assign Pri_elem_10_clock = clock;
  assign Pri_elem_10_reset = reset;
  assign Pri_elem_10_io_pri_update = _T_24 | _T_29; // @[Priority_agent.scala 94:84]
  assign Pri_elem_10_io_pri_update_sig = io_dyn_int_occ_sig; // @[Priority_agent.scala 100:35]
  assign Pri_elem_11_clock = clock;
  assign Pri_elem_11_reset = reset;
  assign Pri_elem_11_io_pri_update = _T_35 | _T_40; // @[Priority_agent.scala 94:84]
  assign Pri_elem_11_io_pri_update_sig = io_dyn_int_occ_sig; // @[Priority_agent.scala 100:35]
  assign Pri_elem_12_clock = clock;
  assign Pri_elem_12_reset = reset;
  assign Pri_elem_12_io_pri_update = _T_46 | _T_51; // @[Priority_agent.scala 94:84]
  assign Pri_elem_12_io_pri_update_sig = io_dyn_int_occ_sig; // @[Priority_agent.scala 100:35]
  assign Pri_elem_13_clock = clock;
  assign Pri_elem_13_reset = reset;
  assign Pri_elem_13_io_pri_update = _T_57 | _T_62; // @[Priority_agent.scala 94:84]
  assign Pri_elem_13_io_pri_update_sig = io_dyn_int_occ_sig; // @[Priority_agent.scala 100:35]
  assign Pri_elem_14_clock = clock;
  assign Pri_elem_14_reset = reset;
  assign Pri_elem_14_io_pri_update = _T_68 | _T_73; // @[Priority_agent.scala 94:84]
  assign Pri_elem_14_io_pri_update_sig = io_dyn_int_occ_sig; // @[Priority_agent.scala 100:35]
  assign Pri_elem_15_clock = clock;
  assign Pri_elem_15_reset = reset;
  assign Pri_elem_15_io_pri_update = _T_79 | _T_84; // @[Priority_agent.scala 94:84]
  assign Pri_elem_15_io_pri_update_sig = io_dyn_int_occ_sig; // @[Priority_agent.scala 100:35]
  assign IntClaimSel_io_ID_in = io_dyn_int_claim_ID; // @[Priority_agent.scala 81:23]
  assign IntOccSel_io_ID_in = io_dyn_int_occ_ID; // @[Priority_agent.scala 80:21]
endmodule
